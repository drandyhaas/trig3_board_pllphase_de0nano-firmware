mux_mhg_inst : mux_mhg PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
